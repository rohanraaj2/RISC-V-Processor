`timescale 1ns / 1ps

`include "Adder.v"
`include "ALU_64_bit.v"
`include "ALU_Control.v"
`include "Branch_module.v"
`include "Control_Unit.v"
`include "Data_Memory.v"
`include "Imm_data_gen.v"
`include "Instruction_Memory.v"
`include "Instruction.v"
`include "MUX.v"
`include "RegisterFile.v"
`include "Program_Counter.v"


module Single_Cycle_Processor(
  
  input clk,
  input reset,
  output reg [63:0] Index_0,
  output reg  [63:0] Index_1,
  output reg  [63:0] Index_2,
  output reg  [63:0] Index_3,
  output reg  [63:0] Index_4,
  output reg  [63:0] Index_5,
  output reg  [63:0] Index_6,
  output reg  [63:0] Index_7,
  output reg  [63:0] Index_8,
  output reg  [63:0] Index_9);
  
  wire [63:0] PC_Out;
  wire [63:0] PC_In;
  wire [63:0] PC_offset_4;
  wire [31:0] IMem_out;
  wire [6:0] opcode;
  wire [4:0] rs1;
  wire [4:0] rs2;
  wire [4:0] rd;
  wire [2:0] funct3;
  wire [6:0] funct7;
  wire [63:0] imm_data;
  wire [1:0] ALUOp;
  wire Branch;
  wire MemRead;
  wire MemtoReg;
  wire MemWrite;
  wire ALUSrc;
  wire RegWrite;
  wire [63:0] write_data;
  wire [63:0] readdata1;
  wire [63:0] readdata2;
  wire [3:0] Operation;
  wire Zero;
  wire [63:0] Result;
  wire [63:0] mux_1_out;
  wire [63:0] DMem_Read;
  wire [63:0] shifted_imm_data;
  wire [63:0] PC_offset_branch;
  wire mux3_select;
  wire bge, blt, bne, beq;
  wire Pos;
  wire [63:0] Index_0;
  wire [63:0] Index_1;
  wire [63:0] Index_2;
  wire [63:0] Index_3;
  wire [63:0] Index_4;
  wire [63:0] Index_5;
  wire [63:0] Index_6;
  wire [63:0] Index_7;
  wire [63:0] Index_8;
  wire [63:0] Index_9;
  wire to_branch;
  
  Adder a1(PC_Out, 64'd4, PC_offset_4);
  MUX m3(PC_offset_4, PC_offset_branch, to_branch, PC_In);
  Program_Counter p1(clk, reset, PC_In, PC_Out);
  Instruction_Memory i1(PC_Out, IMem_out);
  
  Instruction i3(IMem_out, opcode, rd, funct3, rs1, rs2, funct7);
  Imm_data_gen i2(IMem_out, imm_data);
  Control_Unit c1(opcode, ALUOp, Branch, MemRead, MemtoReg, MemWrite, ALUSrc, RegWrite);
  RegisterFile r1(clk, reset, rs1, rs2, rd, write_data, RegWrite, readdata1, readdata2);
  
  Adder a4(PC_Out, imm_data << 1, PC_offset_branch);
  MUX m1(readdata2,	 imm_data, ALUSrc, mux_1_out);

  ALU_Control a2(ALUOp,{IMem_out[30],IMem_out[14:12]},Operation);
  ALU_64_bit a3(readdata1, mux_1_out, Operation, Zero, Result, Pos);
  branch_module b1(Zero, Pos, Branch, funct3, bne, beq, bge, blt, to_branch);

  Data_Memory d1(clk, Result, readdata2, MemWrite, MemRead, DMem_Read, Index_0, Index_1, Index_2, Index_3, Index_4, Index_5, Index_6, Index_7, Index_8, Index_9, funct3);
  MUX m2(Result,DMem_Read,  MemtoReg, write_data);
  
  
endmodule
